`include "register_interface/typedef.svh"
`include "register_interface/assign.svh"

module test_ip_top
    #(
      parameter int unsigned AXI_ADDR_WIDTH = 32,
      localparam int unsigned AXI_DATA_WIDTH = 32,
      parameter int unsigned AXI_ID_WIDTH,
      parameter int unsigned AXI_USER_WIDTH
      )
(
    input clk_i,
    input rst_ni,

    AXI_BUS.Slave axi_slave

);

    import test_ip_reg_pkg::test_ip_reg2hw_t;
    import test_ip_reg_pkg::test_ip_hw2reg_t;

    REG_BUS #(.ADDR_WIDTH(32), .DATA_WIDTH(32)) axi_to_regfile();

    test_ip_reg2hw_t reg_file_to_ip;
    test_ip_hw2reg_t ip_to_reg_file;

    axi_to_reg_intf #(
                      .ADDR_WIDTH(AXI_ADDR_WIDTH),
                      .DATA_WIDTH(AXI_DATA_WIDTH),
                      .ID_WIDTH(AXI_ID_WIDTH),
                      .USER_WIDTH(AXI_USER_WIDTH),
                      .DECOUPLE_W(0)
    ) i_axi2reg (
                 .clk_i,
                 .rst_ni,
                 .testmode_i(test_mode_i),
                 .in(axi_slave),
                 .reg_o(axi_to_regfile)
    );

    //Convert the REG_BUS interface to the struct signals used by autogenerated register file
    typedef logic [AXI_ADDR_WIDTH-1:0] addr_t;
    typedef logic [AXI_DATA_WIDTH-1:0] data_t;
    typedef logic [AXI_DATA_WIDTH/8-1:0] strb_t;
    `REG_BUS_TYPEDEF_REQ(reg_req_t, addr_t, data_t, strb_t);
    `REG_BUS_TYPEDEF_RSP(reg_rsp_t, data_t);
    reg_req_t to_reg_file_req;
    reg_rsp_t from_reg_file_rsp;

    `REG_BUS_ASSIGN_TO_REQ(to_reg_file_req, axi_to_regfile);
    `REG_BUS_ASSIGN_FROM_RSP(axi_to_regfile, from_reg_file_rsp);

    test_ip_reg_top #(
    .reg_req_t(reg_req_t),
    .reg_rsp_t(reg_rsp_t)
    ) i_regfile (
                 .clk_i,
                 .rst_ni,
                 .devmode_i(1'b1),

                 //From the protocol converters to regfile
                 .reg_req_i(to_reg_file_req),
                 .reg_rsp_o(from_reg_file_rsp),

                 //Signals to wide_alu IP
                 .reg2hw(reg_file_to_ip),
                 .hw2reg(ip_to_reg_file)
    );


    test_ip i_test_ip(
        .clk_i,
        .rst_i,
        .reg_a_i(reg_file_to_ip.reg_a.q),
        .reg_b_i(reg_file_to_ip.reg_b.q),
        .res_o(ip_to_reg_file.res.d)
    );
    
endmodule
